//Abdulmalik please do this