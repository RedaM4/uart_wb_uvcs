///Abdulmalik please do this