package uart_module_pkg;

  import uvm_pkg::*;
`include "uvm_macros.svh"


import uart_pkg::*;
import wb_pkg::*;

`include "uart_ver_ref_module.sv"
`include "uart_ver_scoreboard.sv"
`include "uart_ver_ref_env.sv"

endpackage